module adder(input [6:0] I, output [6:0] O);
    assign O = I + 1;
endmodule